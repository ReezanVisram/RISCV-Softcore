`timescale 1ns / 1ps

module data_memory(
    input clk_i,
    input [31:0] address_i,
    input [31:0] data_i,
    output [31:0] data_o
  );

endmodule
