`timescale 1ns / 1ps

module alu(
    input [31:0] data_1_i,
    input [31:0] data_2_i
  );


endmodule
