`timescale 1ns / 1ps

module RISCV_Softcore(
    input clk
  );
  wire [31:0] address;
  wire [31:0] data;



endmodule;
